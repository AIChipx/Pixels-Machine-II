//vector_processor
module vector_processor (a,b);
input a;
output b;
assign b=a;

endmodule 